
task bm_load_test_case1();
    nb = 3;
    nv = 7;
    cmax = 8;
    vmax = 8;

    cbin = '{
        //bin 1
        '{1, 0, 0, 0, 0, 0, 0, 0},
        '{2, 0, 1, 0, 0, 0, 0, 0},
        '{0, 2, 0, 1, 0, 0, 0, 0},
        '{0, 0, 2, 0, 2, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},

        //bin 2
        '{2, 0, 1, 0, 0, 0, 0, 0},
        '{0, 2, 0, 1, 0, 0, 0, 0},
        '{0, 0, 2, 0, 2, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},

        //bin 3
        '{1, 0, 2, 0, 2, 0, 0, 0},
        '{0, 2, 0, 1, 1, 0, 0, 0},
        '{0, 2, 0, 0, 2, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0}
    };

    vbin = '{
        //bin 1
        1, 2, 3, 4, 5, 0, 0, 0,
        //bin 2
        2, 3, 4, 5, 6, 0, 0, 0,
        //bin 3
        1, 2, 5, 6, 7, 0, 0, 0
    };
    run_bm_load();
endtask

