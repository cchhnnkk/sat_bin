
/*** ��������1 ***/

task se_test_case1();

    $display("===============================================");
    $display("test_case 1");

    bin = '{
        '{2, 0, 1, 0, 0, 0, 0, 0},
        '{0, 2, 0, 1, 0, 0, 0, 0},
        '{0, 0, 2, 0, 2, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0}
    };
    //var state list:
    value   = '{0, 0, 0, 0, 0, 0, 0, 0};
    implied = '{0, 0, 0, 0, 0, 0, 0, 0};
    level   = '{0, 0, 0, 0, 0, 0, 0, 0};
    //lvl state list:
    dcd_bin = '{0, 0, 0, 0, 0, 0, 0, 0};
    has_bkt = '{0, 0, 0, 0, 0, 0, 0, 0};
    //ctrl
    cur_bin_num = 1;
    load_lvl = 1;
    base_lvl = 1;

    //�����������
    process_len = 6;
    process_data = '{
        '{"decision", 0, 1, 2},
        '{"bcp",      2, 1, 2},
        '{"bcp",      4, 2, 2},
        '{"decision", 1, 1, 3},
        '{"bcp",      3, 1, 3},
        '{"psat",     0, 0, 0}
    };

    run_test_case();
endtask
