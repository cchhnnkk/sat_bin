
/*** 测试数据7 ***/

task se_test_case7();

    $display("===============================================");
    $display("test_case 7");

	bin = '{
		'{0, 1, 0, 1, 0, 0, 1, 0},
		'{0, 2, 1, 0, 1, 0, 0, 0},
		'{1, 0, 2, 0, 0, 2, 0, 0},
		'{0, 0, 0, 0, 0, 0, 0, 0},
		'{0, 0, 0, 0, 0, 0, 0, 0},
		'{0, 0, 0, 0, 0, 0, 0, 0},
		'{0, 0, 0, 0, 0, 0, 0, 0},
		'{0, 0, 0, 0, 0, 0, 0, 0}
	};
	//var state list:
	value   = '{2, 1, 0, 2, 0, 1, 1, 0};
	implied = '{0, 0, 0, 1, 0, 1, 1, 0};
	level   = '{4, 2, 0, 3, 0, 5, 5, 0};
	//lvl state list:
	dcd_bin = '{7, 10, 11, 14, 14, 0, 0, 0};
	has_bkt = '{1, 1, 1, 1, 0, 0, 0, 0};
	//ctrl
	cur_bin_num = 23;
	base_lvl = 8;
	load_lvl = 8;

    //运算过程数据
    process_len = 3;
    process_data = '{
        '{"bcp",      2, 2, 5},
        '{"bcp",      1, 1, 5},
        '{"psat",     0, 0, 0}
    };

    run_test_case();
endtask

